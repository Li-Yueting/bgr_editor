magic
tech sky130A
magscale 1 2
timestamp 1656304247
<< nwell >>
rect 120 1707 3094 1940
rect 120 294 3095 1707
rect 217 293 3095 294
<< pmoslvt >>
rect 311 355 711 1645
rect 769 355 1169 1645
rect 1227 355 1627 1645
rect 1685 355 2085 1645
rect 2143 355 2543 1645
rect 2601 355 3001 1645
<< pdiff >>
rect 253 1629 311 1645
rect 253 1595 265 1629
rect 299 1595 311 1629
rect 253 1561 311 1595
rect 253 1527 265 1561
rect 299 1527 311 1561
rect 253 1493 311 1527
rect 253 1459 265 1493
rect 299 1459 311 1493
rect 253 1425 311 1459
rect 253 1391 265 1425
rect 299 1391 311 1425
rect 253 1357 311 1391
rect 253 1323 265 1357
rect 299 1323 311 1357
rect 253 1289 311 1323
rect 253 1255 265 1289
rect 299 1255 311 1289
rect 253 1221 311 1255
rect 253 1187 265 1221
rect 299 1187 311 1221
rect 253 1153 311 1187
rect 253 1119 265 1153
rect 299 1119 311 1153
rect 253 1085 311 1119
rect 253 1051 265 1085
rect 299 1051 311 1085
rect 253 1017 311 1051
rect 253 983 265 1017
rect 299 983 311 1017
rect 253 949 311 983
rect 253 915 265 949
rect 299 915 311 949
rect 253 881 311 915
rect 253 847 265 881
rect 299 847 311 881
rect 253 813 311 847
rect 253 779 265 813
rect 299 779 311 813
rect 253 745 311 779
rect 253 711 265 745
rect 299 711 311 745
rect 253 677 311 711
rect 253 643 265 677
rect 299 643 311 677
rect 253 609 311 643
rect 253 575 265 609
rect 299 575 311 609
rect 253 541 311 575
rect 253 507 265 541
rect 299 507 311 541
rect 253 473 311 507
rect 253 439 265 473
rect 299 439 311 473
rect 253 405 311 439
rect 253 371 265 405
rect 299 371 311 405
rect 253 355 311 371
rect 711 1629 769 1645
rect 711 1595 723 1629
rect 757 1595 769 1629
rect 711 1561 769 1595
rect 711 1527 723 1561
rect 757 1527 769 1561
rect 711 1493 769 1527
rect 711 1459 723 1493
rect 757 1459 769 1493
rect 711 1425 769 1459
rect 711 1391 723 1425
rect 757 1391 769 1425
rect 711 1357 769 1391
rect 711 1323 723 1357
rect 757 1323 769 1357
rect 711 1289 769 1323
rect 711 1255 723 1289
rect 757 1255 769 1289
rect 711 1221 769 1255
rect 711 1187 723 1221
rect 757 1187 769 1221
rect 711 1153 769 1187
rect 711 1119 723 1153
rect 757 1119 769 1153
rect 711 1085 769 1119
rect 711 1051 723 1085
rect 757 1051 769 1085
rect 711 1017 769 1051
rect 711 983 723 1017
rect 757 983 769 1017
rect 711 949 769 983
rect 711 915 723 949
rect 757 915 769 949
rect 711 881 769 915
rect 711 847 723 881
rect 757 847 769 881
rect 711 813 769 847
rect 711 779 723 813
rect 757 779 769 813
rect 711 745 769 779
rect 711 711 723 745
rect 757 711 769 745
rect 711 677 769 711
rect 711 643 723 677
rect 757 643 769 677
rect 711 609 769 643
rect 711 575 723 609
rect 757 575 769 609
rect 711 541 769 575
rect 711 507 723 541
rect 757 507 769 541
rect 711 473 769 507
rect 711 439 723 473
rect 757 439 769 473
rect 711 405 769 439
rect 711 371 723 405
rect 757 371 769 405
rect 711 355 769 371
rect 1169 1629 1227 1645
rect 1169 1595 1181 1629
rect 1215 1595 1227 1629
rect 1169 1561 1227 1595
rect 1169 1527 1181 1561
rect 1215 1527 1227 1561
rect 1169 1493 1227 1527
rect 1169 1459 1181 1493
rect 1215 1459 1227 1493
rect 1169 1425 1227 1459
rect 1169 1391 1181 1425
rect 1215 1391 1227 1425
rect 1169 1357 1227 1391
rect 1169 1323 1181 1357
rect 1215 1323 1227 1357
rect 1169 1289 1227 1323
rect 1169 1255 1181 1289
rect 1215 1255 1227 1289
rect 1169 1221 1227 1255
rect 1169 1187 1181 1221
rect 1215 1187 1227 1221
rect 1169 1153 1227 1187
rect 1169 1119 1181 1153
rect 1215 1119 1227 1153
rect 1169 1085 1227 1119
rect 1169 1051 1181 1085
rect 1215 1051 1227 1085
rect 1169 1017 1227 1051
rect 1169 983 1181 1017
rect 1215 983 1227 1017
rect 1169 949 1227 983
rect 1169 915 1181 949
rect 1215 915 1227 949
rect 1169 881 1227 915
rect 1169 847 1181 881
rect 1215 847 1227 881
rect 1169 813 1227 847
rect 1169 779 1181 813
rect 1215 779 1227 813
rect 1169 745 1227 779
rect 1169 711 1181 745
rect 1215 711 1227 745
rect 1169 677 1227 711
rect 1169 643 1181 677
rect 1215 643 1227 677
rect 1169 609 1227 643
rect 1169 575 1181 609
rect 1215 575 1227 609
rect 1169 541 1227 575
rect 1169 507 1181 541
rect 1215 507 1227 541
rect 1169 473 1227 507
rect 1169 439 1181 473
rect 1215 439 1227 473
rect 1169 405 1227 439
rect 1169 371 1181 405
rect 1215 371 1227 405
rect 1169 355 1227 371
rect 1627 1629 1685 1645
rect 1627 1595 1639 1629
rect 1673 1595 1685 1629
rect 1627 1561 1685 1595
rect 1627 1527 1639 1561
rect 1673 1527 1685 1561
rect 1627 1493 1685 1527
rect 1627 1459 1639 1493
rect 1673 1459 1685 1493
rect 1627 1425 1685 1459
rect 1627 1391 1639 1425
rect 1673 1391 1685 1425
rect 1627 1357 1685 1391
rect 1627 1323 1639 1357
rect 1673 1323 1685 1357
rect 1627 1289 1685 1323
rect 1627 1255 1639 1289
rect 1673 1255 1685 1289
rect 1627 1221 1685 1255
rect 1627 1187 1639 1221
rect 1673 1187 1685 1221
rect 1627 1153 1685 1187
rect 1627 1119 1639 1153
rect 1673 1119 1685 1153
rect 1627 1085 1685 1119
rect 1627 1051 1639 1085
rect 1673 1051 1685 1085
rect 1627 1017 1685 1051
rect 1627 983 1639 1017
rect 1673 983 1685 1017
rect 1627 949 1685 983
rect 1627 915 1639 949
rect 1673 915 1685 949
rect 1627 881 1685 915
rect 1627 847 1639 881
rect 1673 847 1685 881
rect 1627 813 1685 847
rect 1627 779 1639 813
rect 1673 779 1685 813
rect 1627 745 1685 779
rect 1627 711 1639 745
rect 1673 711 1685 745
rect 1627 677 1685 711
rect 1627 643 1639 677
rect 1673 643 1685 677
rect 1627 609 1685 643
rect 1627 575 1639 609
rect 1673 575 1685 609
rect 1627 541 1685 575
rect 1627 507 1639 541
rect 1673 507 1685 541
rect 1627 473 1685 507
rect 1627 439 1639 473
rect 1673 439 1685 473
rect 1627 405 1685 439
rect 1627 371 1639 405
rect 1673 371 1685 405
rect 1627 355 1685 371
rect 2085 1629 2143 1645
rect 2085 1595 2097 1629
rect 2131 1595 2143 1629
rect 2085 1561 2143 1595
rect 2085 1527 2097 1561
rect 2131 1527 2143 1561
rect 2085 1493 2143 1527
rect 2085 1459 2097 1493
rect 2131 1459 2143 1493
rect 2085 1425 2143 1459
rect 2085 1391 2097 1425
rect 2131 1391 2143 1425
rect 2085 1357 2143 1391
rect 2085 1323 2097 1357
rect 2131 1323 2143 1357
rect 2085 1289 2143 1323
rect 2085 1255 2097 1289
rect 2131 1255 2143 1289
rect 2085 1221 2143 1255
rect 2085 1187 2097 1221
rect 2131 1187 2143 1221
rect 2085 1153 2143 1187
rect 2085 1119 2097 1153
rect 2131 1119 2143 1153
rect 2085 1085 2143 1119
rect 2085 1051 2097 1085
rect 2131 1051 2143 1085
rect 2085 1017 2143 1051
rect 2085 983 2097 1017
rect 2131 983 2143 1017
rect 2085 949 2143 983
rect 2085 915 2097 949
rect 2131 915 2143 949
rect 2085 881 2143 915
rect 2085 847 2097 881
rect 2131 847 2143 881
rect 2085 813 2143 847
rect 2085 779 2097 813
rect 2131 779 2143 813
rect 2085 745 2143 779
rect 2085 711 2097 745
rect 2131 711 2143 745
rect 2085 677 2143 711
rect 2085 643 2097 677
rect 2131 643 2143 677
rect 2085 609 2143 643
rect 2085 575 2097 609
rect 2131 575 2143 609
rect 2085 541 2143 575
rect 2085 507 2097 541
rect 2131 507 2143 541
rect 2085 473 2143 507
rect 2085 439 2097 473
rect 2131 439 2143 473
rect 2085 405 2143 439
rect 2085 371 2097 405
rect 2131 371 2143 405
rect 2085 355 2143 371
rect 2543 1629 2601 1645
rect 2543 1595 2555 1629
rect 2589 1595 2601 1629
rect 2543 1561 2601 1595
rect 2543 1527 2555 1561
rect 2589 1527 2601 1561
rect 2543 1493 2601 1527
rect 2543 1459 2555 1493
rect 2589 1459 2601 1493
rect 2543 1425 2601 1459
rect 2543 1391 2555 1425
rect 2589 1391 2601 1425
rect 2543 1357 2601 1391
rect 2543 1323 2555 1357
rect 2589 1323 2601 1357
rect 2543 1289 2601 1323
rect 2543 1255 2555 1289
rect 2589 1255 2601 1289
rect 2543 1221 2601 1255
rect 2543 1187 2555 1221
rect 2589 1187 2601 1221
rect 2543 1153 2601 1187
rect 2543 1119 2555 1153
rect 2589 1119 2601 1153
rect 2543 1085 2601 1119
rect 2543 1051 2555 1085
rect 2589 1051 2601 1085
rect 2543 1017 2601 1051
rect 2543 983 2555 1017
rect 2589 983 2601 1017
rect 2543 949 2601 983
rect 2543 915 2555 949
rect 2589 915 2601 949
rect 2543 881 2601 915
rect 2543 847 2555 881
rect 2589 847 2601 881
rect 2543 813 2601 847
rect 2543 779 2555 813
rect 2589 779 2601 813
rect 2543 745 2601 779
rect 2543 711 2555 745
rect 2589 711 2601 745
rect 2543 677 2601 711
rect 2543 643 2555 677
rect 2589 643 2601 677
rect 2543 609 2601 643
rect 2543 575 2555 609
rect 2589 575 2601 609
rect 2543 541 2601 575
rect 2543 507 2555 541
rect 2589 507 2601 541
rect 2543 473 2601 507
rect 2543 439 2555 473
rect 2589 439 2601 473
rect 2543 405 2601 439
rect 2543 371 2555 405
rect 2589 371 2601 405
rect 2543 355 2601 371
rect 3001 1629 3059 1645
rect 3001 1595 3013 1629
rect 3047 1595 3059 1629
rect 3001 1561 3059 1595
rect 3001 1527 3013 1561
rect 3047 1527 3059 1561
rect 3001 1493 3059 1527
rect 3001 1459 3013 1493
rect 3047 1459 3059 1493
rect 3001 1425 3059 1459
rect 3001 1391 3013 1425
rect 3047 1391 3059 1425
rect 3001 1357 3059 1391
rect 3001 1323 3013 1357
rect 3047 1323 3059 1357
rect 3001 1289 3059 1323
rect 3001 1255 3013 1289
rect 3047 1255 3059 1289
rect 3001 1221 3059 1255
rect 3001 1187 3013 1221
rect 3047 1187 3059 1221
rect 3001 1153 3059 1187
rect 3001 1119 3013 1153
rect 3047 1119 3059 1153
rect 3001 1085 3059 1119
rect 3001 1051 3013 1085
rect 3047 1051 3059 1085
rect 3001 1017 3059 1051
rect 3001 983 3013 1017
rect 3047 983 3059 1017
rect 3001 949 3059 983
rect 3001 915 3013 949
rect 3047 915 3059 949
rect 3001 881 3059 915
rect 3001 847 3013 881
rect 3047 847 3059 881
rect 3001 813 3059 847
rect 3001 779 3013 813
rect 3047 779 3059 813
rect 3001 745 3059 779
rect 3001 711 3013 745
rect 3047 711 3059 745
rect 3001 677 3059 711
rect 3001 643 3013 677
rect 3047 643 3059 677
rect 3001 609 3059 643
rect 3001 575 3013 609
rect 3047 575 3059 609
rect 3001 541 3059 575
rect 3001 507 3013 541
rect 3047 507 3059 541
rect 3001 473 3059 507
rect 3001 439 3013 473
rect 3047 439 3059 473
rect 3001 405 3059 439
rect 3001 371 3013 405
rect 3047 371 3059 405
rect 3001 355 3059 371
<< pdiffc >>
rect 265 1595 299 1629
rect 265 1527 299 1561
rect 265 1459 299 1493
rect 265 1391 299 1425
rect 265 1323 299 1357
rect 265 1255 299 1289
rect 265 1187 299 1221
rect 265 1119 299 1153
rect 265 1051 299 1085
rect 265 983 299 1017
rect 265 915 299 949
rect 265 847 299 881
rect 265 779 299 813
rect 265 711 299 745
rect 265 643 299 677
rect 265 575 299 609
rect 265 507 299 541
rect 265 439 299 473
rect 265 371 299 405
rect 723 1595 757 1629
rect 723 1527 757 1561
rect 723 1459 757 1493
rect 723 1391 757 1425
rect 723 1323 757 1357
rect 723 1255 757 1289
rect 723 1187 757 1221
rect 723 1119 757 1153
rect 723 1051 757 1085
rect 723 983 757 1017
rect 723 915 757 949
rect 723 847 757 881
rect 723 779 757 813
rect 723 711 757 745
rect 723 643 757 677
rect 723 575 757 609
rect 723 507 757 541
rect 723 439 757 473
rect 723 371 757 405
rect 1181 1595 1215 1629
rect 1181 1527 1215 1561
rect 1181 1459 1215 1493
rect 1181 1391 1215 1425
rect 1181 1323 1215 1357
rect 1181 1255 1215 1289
rect 1181 1187 1215 1221
rect 1181 1119 1215 1153
rect 1181 1051 1215 1085
rect 1181 983 1215 1017
rect 1181 915 1215 949
rect 1181 847 1215 881
rect 1181 779 1215 813
rect 1181 711 1215 745
rect 1181 643 1215 677
rect 1181 575 1215 609
rect 1181 507 1215 541
rect 1181 439 1215 473
rect 1181 371 1215 405
rect 1639 1595 1673 1629
rect 1639 1527 1673 1561
rect 1639 1459 1673 1493
rect 1639 1391 1673 1425
rect 1639 1323 1673 1357
rect 1639 1255 1673 1289
rect 1639 1187 1673 1221
rect 1639 1119 1673 1153
rect 1639 1051 1673 1085
rect 1639 983 1673 1017
rect 1639 915 1673 949
rect 1639 847 1673 881
rect 1639 779 1673 813
rect 1639 711 1673 745
rect 1639 643 1673 677
rect 1639 575 1673 609
rect 1639 507 1673 541
rect 1639 439 1673 473
rect 1639 371 1673 405
rect 2097 1595 2131 1629
rect 2097 1527 2131 1561
rect 2097 1459 2131 1493
rect 2097 1391 2131 1425
rect 2097 1323 2131 1357
rect 2097 1255 2131 1289
rect 2097 1187 2131 1221
rect 2097 1119 2131 1153
rect 2097 1051 2131 1085
rect 2097 983 2131 1017
rect 2097 915 2131 949
rect 2097 847 2131 881
rect 2097 779 2131 813
rect 2097 711 2131 745
rect 2097 643 2131 677
rect 2097 575 2131 609
rect 2097 507 2131 541
rect 2097 439 2131 473
rect 2097 371 2131 405
rect 2555 1595 2589 1629
rect 2555 1527 2589 1561
rect 2555 1459 2589 1493
rect 2555 1391 2589 1425
rect 2555 1323 2589 1357
rect 2555 1255 2589 1289
rect 2555 1187 2589 1221
rect 2555 1119 2589 1153
rect 2555 1051 2589 1085
rect 2555 983 2589 1017
rect 2555 915 2589 949
rect 2555 847 2589 881
rect 2555 779 2589 813
rect 2555 711 2589 745
rect 2555 643 2589 677
rect 2555 575 2589 609
rect 2555 507 2589 541
rect 2555 439 2589 473
rect 2555 371 2589 405
rect 3013 1595 3047 1629
rect 3013 1527 3047 1561
rect 3013 1459 3047 1493
rect 3013 1391 3047 1425
rect 3013 1323 3047 1357
rect 3013 1255 3047 1289
rect 3013 1187 3047 1221
rect 3013 1119 3047 1153
rect 3013 1051 3047 1085
rect 3013 983 3047 1017
rect 3013 915 3047 949
rect 3013 847 3047 881
rect 3013 779 3047 813
rect 3013 711 3047 745
rect 3013 643 3047 677
rect 3013 575 3047 609
rect 3013 507 3047 541
rect 3013 439 3047 473
rect 3013 371 3047 405
<< nsubdiff >>
rect 1216 1807 1336 1810
rect 158 1757 198 1800
rect 1216 1773 1261 1807
rect 1295 1773 1336 1807
rect 1216 1770 1336 1773
rect 158 1723 161 1757
rect 195 1723 198 1757
rect 158 1680 198 1723
<< nsubdiffcont >>
rect 1261 1773 1295 1807
rect 161 1723 195 1757
<< poly >>
rect 311 1645 711 1671
rect 769 1645 1169 1671
rect 1227 1645 1627 1671
rect 1685 1645 2085 1671
rect 2143 1645 2543 1671
rect 2601 1645 3001 1671
rect 311 329 711 355
rect 769 329 1169 355
rect 1227 329 1627 355
rect 1685 329 2085 355
rect 2143 329 2543 355
rect 2601 329 3001 355
rect 458 184 578 329
rect 914 184 1034 329
rect 1370 184 1490 329
rect 1826 184 1946 329
rect 2282 184 2402 329
rect 2738 184 2858 329
rect 218 151 3094 184
rect 218 117 401 151
rect 435 117 801 151
rect 835 117 1201 151
rect 1235 117 1601 151
rect 1635 117 2001 151
rect 2035 117 2401 151
rect 2435 117 2801 151
rect 2835 117 3094 151
rect 218 84 3094 117
<< polycont >>
rect 401 117 435 151
rect 801 117 835 151
rect 1201 117 1235 151
rect 1601 117 1635 151
rect 2001 117 2035 151
rect 2401 117 2435 151
rect 2801 117 2835 151
<< locali >>
rect 120 1897 3094 1910
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3094 1897
rect 120 1850 3094 1863
rect 148 1757 208 1850
rect 1196 1807 1356 1850
rect 1196 1773 1261 1807
rect 1295 1773 1356 1807
rect 1196 1770 1356 1773
rect 148 1723 161 1757
rect 195 1723 208 1757
rect 148 1640 208 1723
rect 278 1690 3094 1730
rect 265 1629 299 1649
rect 265 1561 299 1595
rect 265 1493 299 1523
rect 265 1425 299 1451
rect 265 1357 299 1379
rect 265 1289 299 1307
rect 265 1221 299 1235
rect 265 1153 299 1163
rect 265 1085 299 1091
rect 265 1017 299 1019
rect 265 981 299 983
rect 265 909 299 915
rect 265 837 299 847
rect 265 765 299 779
rect 265 693 299 711
rect 265 621 299 643
rect 265 549 299 575
rect 265 477 299 507
rect 265 405 299 439
rect 265 270 299 371
rect 723 1629 757 1690
rect 723 1561 757 1595
rect 723 1493 757 1523
rect 723 1425 757 1451
rect 723 1357 757 1379
rect 723 1289 757 1307
rect 723 1221 757 1235
rect 723 1153 757 1163
rect 723 1085 757 1091
rect 723 1017 757 1019
rect 723 981 757 983
rect 723 909 757 915
rect 723 837 757 847
rect 723 765 757 779
rect 723 693 757 711
rect 723 621 757 643
rect 723 549 757 575
rect 723 477 757 507
rect 723 405 757 439
rect 723 351 757 371
rect 1181 1629 1215 1649
rect 1181 1561 1215 1595
rect 1181 1493 1215 1523
rect 1181 1425 1215 1451
rect 1181 1357 1215 1379
rect 1181 1289 1215 1307
rect 1181 1221 1215 1235
rect 1181 1153 1215 1163
rect 1181 1085 1215 1091
rect 1181 1017 1215 1019
rect 1181 981 1215 983
rect 1181 909 1215 915
rect 1181 837 1215 847
rect 1181 765 1215 779
rect 1181 693 1215 711
rect 1181 621 1215 643
rect 1181 549 1215 575
rect 1181 477 1215 507
rect 1181 405 1215 439
rect 1181 270 1215 371
rect 1639 1629 1673 1690
rect 1639 1561 1673 1595
rect 1639 1493 1673 1523
rect 1639 1425 1673 1451
rect 1639 1357 1673 1379
rect 1639 1289 1673 1307
rect 1639 1221 1673 1235
rect 1639 1153 1673 1163
rect 1639 1085 1673 1091
rect 1639 1017 1673 1019
rect 1639 981 1673 983
rect 1639 909 1673 915
rect 1639 837 1673 847
rect 1639 765 1673 779
rect 1639 693 1673 711
rect 1639 621 1673 643
rect 1639 549 1673 575
rect 1639 477 1673 507
rect 1639 405 1673 439
rect 1639 351 1673 371
rect 2097 1629 2131 1649
rect 2097 1561 2131 1595
rect 2097 1493 2131 1523
rect 2097 1425 2131 1451
rect 2097 1357 2131 1379
rect 2097 1289 2131 1307
rect 2097 1221 2131 1235
rect 2097 1153 2131 1163
rect 2097 1085 2131 1091
rect 2097 1017 2131 1019
rect 2097 981 2131 983
rect 2097 909 2131 915
rect 2097 837 2131 847
rect 2097 765 2131 779
rect 2097 693 2131 711
rect 2097 621 2131 643
rect 2097 549 2131 575
rect 2097 477 2131 507
rect 2097 405 2131 439
rect 2097 270 2131 371
rect 2555 1629 2589 1690
rect 2555 1561 2589 1595
rect 2555 1493 2589 1523
rect 2555 1425 2589 1451
rect 2555 1357 2589 1379
rect 2555 1289 2589 1307
rect 2555 1221 2589 1235
rect 2555 1153 2589 1163
rect 2555 1085 2589 1091
rect 2555 1017 2589 1019
rect 2555 981 2589 983
rect 2555 909 2589 915
rect 2555 837 2589 847
rect 2555 765 2589 779
rect 2555 693 2589 711
rect 2555 621 2589 643
rect 2555 549 2589 575
rect 2555 477 2589 507
rect 2555 405 2589 439
rect 2555 351 2589 371
rect 3013 1629 3047 1649
rect 3013 1561 3047 1595
rect 3013 1493 3047 1523
rect 3013 1425 3047 1451
rect 3013 1357 3047 1379
rect 3013 1289 3047 1307
rect 3013 1221 3047 1235
rect 3013 1153 3047 1163
rect 3013 1085 3047 1091
rect 3013 1017 3047 1019
rect 3013 981 3047 983
rect 3013 909 3047 915
rect 3013 837 3047 847
rect 3013 765 3047 779
rect 3013 693 3047 711
rect 3013 621 3047 643
rect 3013 549 3047 575
rect 3013 477 3047 507
rect 3013 405 3047 439
rect 3013 270 3047 371
rect 218 210 3094 270
rect 218 151 3094 164
rect 218 117 401 151
rect 435 117 801 151
rect 835 117 1201 151
rect 1235 117 1601 151
rect 1635 117 2001 151
rect 2035 117 2401 151
rect 2435 117 2801 151
rect 2835 117 3094 151
rect 218 104 3094 117
rect 120 17 3094 30
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3094 17
rect 120 -30 3094 -17
<< viali >>
rect 401 1863 435 1897
rect 801 1863 835 1897
rect 1201 1863 1235 1897
rect 1601 1863 1635 1897
rect 2001 1863 2035 1897
rect 2401 1863 2435 1897
rect 2801 1863 2835 1897
rect 265 1595 299 1629
rect 265 1527 299 1557
rect 265 1523 299 1527
rect 265 1459 299 1485
rect 265 1451 299 1459
rect 265 1391 299 1413
rect 265 1379 299 1391
rect 265 1323 299 1341
rect 265 1307 299 1323
rect 265 1255 299 1269
rect 265 1235 299 1255
rect 265 1187 299 1197
rect 265 1163 299 1187
rect 265 1119 299 1125
rect 265 1091 299 1119
rect 265 1051 299 1053
rect 265 1019 299 1051
rect 265 949 299 981
rect 265 947 299 949
rect 265 881 299 909
rect 265 875 299 881
rect 265 813 299 837
rect 265 803 299 813
rect 265 745 299 765
rect 265 731 299 745
rect 265 677 299 693
rect 265 659 299 677
rect 265 609 299 621
rect 265 587 299 609
rect 265 541 299 549
rect 265 515 299 541
rect 265 473 299 477
rect 265 443 299 473
rect 265 371 299 405
rect 723 1595 757 1629
rect 723 1527 757 1557
rect 723 1523 757 1527
rect 723 1459 757 1485
rect 723 1451 757 1459
rect 723 1391 757 1413
rect 723 1379 757 1391
rect 723 1323 757 1341
rect 723 1307 757 1323
rect 723 1255 757 1269
rect 723 1235 757 1255
rect 723 1187 757 1197
rect 723 1163 757 1187
rect 723 1119 757 1125
rect 723 1091 757 1119
rect 723 1051 757 1053
rect 723 1019 757 1051
rect 723 949 757 981
rect 723 947 757 949
rect 723 881 757 909
rect 723 875 757 881
rect 723 813 757 837
rect 723 803 757 813
rect 723 745 757 765
rect 723 731 757 745
rect 723 677 757 693
rect 723 659 757 677
rect 723 609 757 621
rect 723 587 757 609
rect 723 541 757 549
rect 723 515 757 541
rect 723 473 757 477
rect 723 443 757 473
rect 723 371 757 405
rect 1181 1595 1215 1629
rect 1181 1527 1215 1557
rect 1181 1523 1215 1527
rect 1181 1459 1215 1485
rect 1181 1451 1215 1459
rect 1181 1391 1215 1413
rect 1181 1379 1215 1391
rect 1181 1323 1215 1341
rect 1181 1307 1215 1323
rect 1181 1255 1215 1269
rect 1181 1235 1215 1255
rect 1181 1187 1215 1197
rect 1181 1163 1215 1187
rect 1181 1119 1215 1125
rect 1181 1091 1215 1119
rect 1181 1051 1215 1053
rect 1181 1019 1215 1051
rect 1181 949 1215 981
rect 1181 947 1215 949
rect 1181 881 1215 909
rect 1181 875 1215 881
rect 1181 813 1215 837
rect 1181 803 1215 813
rect 1181 745 1215 765
rect 1181 731 1215 745
rect 1181 677 1215 693
rect 1181 659 1215 677
rect 1181 609 1215 621
rect 1181 587 1215 609
rect 1181 541 1215 549
rect 1181 515 1215 541
rect 1181 473 1215 477
rect 1181 443 1215 473
rect 1181 371 1215 405
rect 1639 1595 1673 1629
rect 1639 1527 1673 1557
rect 1639 1523 1673 1527
rect 1639 1459 1673 1485
rect 1639 1451 1673 1459
rect 1639 1391 1673 1413
rect 1639 1379 1673 1391
rect 1639 1323 1673 1341
rect 1639 1307 1673 1323
rect 1639 1255 1673 1269
rect 1639 1235 1673 1255
rect 1639 1187 1673 1197
rect 1639 1163 1673 1187
rect 1639 1119 1673 1125
rect 1639 1091 1673 1119
rect 1639 1051 1673 1053
rect 1639 1019 1673 1051
rect 1639 949 1673 981
rect 1639 947 1673 949
rect 1639 881 1673 909
rect 1639 875 1673 881
rect 1639 813 1673 837
rect 1639 803 1673 813
rect 1639 745 1673 765
rect 1639 731 1673 745
rect 1639 677 1673 693
rect 1639 659 1673 677
rect 1639 609 1673 621
rect 1639 587 1673 609
rect 1639 541 1673 549
rect 1639 515 1673 541
rect 1639 473 1673 477
rect 1639 443 1673 473
rect 1639 371 1673 405
rect 2097 1595 2131 1629
rect 2097 1527 2131 1557
rect 2097 1523 2131 1527
rect 2097 1459 2131 1485
rect 2097 1451 2131 1459
rect 2097 1391 2131 1413
rect 2097 1379 2131 1391
rect 2097 1323 2131 1341
rect 2097 1307 2131 1323
rect 2097 1255 2131 1269
rect 2097 1235 2131 1255
rect 2097 1187 2131 1197
rect 2097 1163 2131 1187
rect 2097 1119 2131 1125
rect 2097 1091 2131 1119
rect 2097 1051 2131 1053
rect 2097 1019 2131 1051
rect 2097 949 2131 981
rect 2097 947 2131 949
rect 2097 881 2131 909
rect 2097 875 2131 881
rect 2097 813 2131 837
rect 2097 803 2131 813
rect 2097 745 2131 765
rect 2097 731 2131 745
rect 2097 677 2131 693
rect 2097 659 2131 677
rect 2097 609 2131 621
rect 2097 587 2131 609
rect 2097 541 2131 549
rect 2097 515 2131 541
rect 2097 473 2131 477
rect 2097 443 2131 473
rect 2097 371 2131 405
rect 2555 1595 2589 1629
rect 2555 1527 2589 1557
rect 2555 1523 2589 1527
rect 2555 1459 2589 1485
rect 2555 1451 2589 1459
rect 2555 1391 2589 1413
rect 2555 1379 2589 1391
rect 2555 1323 2589 1341
rect 2555 1307 2589 1323
rect 2555 1255 2589 1269
rect 2555 1235 2589 1255
rect 2555 1187 2589 1197
rect 2555 1163 2589 1187
rect 2555 1119 2589 1125
rect 2555 1091 2589 1119
rect 2555 1051 2589 1053
rect 2555 1019 2589 1051
rect 2555 949 2589 981
rect 2555 947 2589 949
rect 2555 881 2589 909
rect 2555 875 2589 881
rect 2555 813 2589 837
rect 2555 803 2589 813
rect 2555 745 2589 765
rect 2555 731 2589 745
rect 2555 677 2589 693
rect 2555 659 2589 677
rect 2555 609 2589 621
rect 2555 587 2589 609
rect 2555 541 2589 549
rect 2555 515 2589 541
rect 2555 473 2589 477
rect 2555 443 2589 473
rect 2555 371 2589 405
rect 3013 1595 3047 1629
rect 3013 1527 3047 1557
rect 3013 1523 3047 1527
rect 3013 1459 3047 1485
rect 3013 1451 3047 1459
rect 3013 1391 3047 1413
rect 3013 1379 3047 1391
rect 3013 1323 3047 1341
rect 3013 1307 3047 1323
rect 3013 1255 3047 1269
rect 3013 1235 3047 1255
rect 3013 1187 3047 1197
rect 3013 1163 3047 1187
rect 3013 1119 3047 1125
rect 3013 1091 3047 1119
rect 3013 1051 3047 1053
rect 3013 1019 3047 1051
rect 3013 949 3047 981
rect 3013 947 3047 949
rect 3013 881 3047 909
rect 3013 875 3047 881
rect 3013 813 3047 837
rect 3013 803 3047 813
rect 3013 745 3047 765
rect 3013 731 3047 745
rect 3013 677 3047 693
rect 3013 659 3047 677
rect 3013 609 3047 621
rect 3013 587 3047 609
rect 3013 541 3047 549
rect 3013 515 3047 541
rect 3013 473 3047 477
rect 3013 443 3047 473
rect 3013 371 3047 405
rect 401 -17 435 17
rect 801 -17 835 17
rect 1201 -17 1235 17
rect 1601 -17 1635 17
rect 2001 -17 2035 17
rect 2401 -17 2435 17
rect 2801 -17 2835 17
<< metal1 >>
rect 120 1897 3094 1940
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3094 1897
rect 120 1820 3094 1863
rect 259 1629 305 1645
rect 259 1595 265 1629
rect 299 1595 305 1629
rect 259 1557 305 1595
rect 259 1523 265 1557
rect 299 1523 305 1557
rect 259 1485 305 1523
rect 259 1451 265 1485
rect 299 1451 305 1485
rect 259 1413 305 1451
rect 259 1379 265 1413
rect 299 1379 305 1413
rect 259 1341 305 1379
rect 259 1307 265 1341
rect 299 1307 305 1341
rect 259 1269 305 1307
rect 259 1235 265 1269
rect 299 1235 305 1269
rect 259 1197 305 1235
rect 259 1163 265 1197
rect 299 1163 305 1197
rect 259 1125 305 1163
rect 259 1091 265 1125
rect 299 1091 305 1125
rect 259 1053 305 1091
rect 259 1019 265 1053
rect 299 1019 305 1053
rect 259 981 305 1019
rect 259 947 265 981
rect 299 947 305 981
rect 259 909 305 947
rect 259 875 265 909
rect 299 875 305 909
rect 259 837 305 875
rect 259 803 265 837
rect 299 803 305 837
rect 259 765 305 803
rect 259 731 265 765
rect 299 731 305 765
rect 259 693 305 731
rect 259 659 265 693
rect 299 659 305 693
rect 259 621 305 659
rect 259 587 265 621
rect 299 587 305 621
rect 259 549 305 587
rect 259 515 265 549
rect 299 515 305 549
rect 259 477 305 515
rect 259 443 265 477
rect 299 443 305 477
rect 259 405 305 443
rect 259 371 265 405
rect 299 371 305 405
rect 259 355 305 371
rect 717 1629 763 1645
rect 717 1595 723 1629
rect 757 1595 763 1629
rect 717 1557 763 1595
rect 717 1523 723 1557
rect 757 1523 763 1557
rect 717 1485 763 1523
rect 717 1451 723 1485
rect 757 1451 763 1485
rect 717 1413 763 1451
rect 717 1379 723 1413
rect 757 1379 763 1413
rect 717 1341 763 1379
rect 717 1307 723 1341
rect 757 1307 763 1341
rect 717 1269 763 1307
rect 717 1235 723 1269
rect 757 1235 763 1269
rect 717 1197 763 1235
rect 717 1163 723 1197
rect 757 1163 763 1197
rect 717 1125 763 1163
rect 717 1091 723 1125
rect 757 1091 763 1125
rect 717 1053 763 1091
rect 717 1019 723 1053
rect 757 1019 763 1053
rect 717 981 763 1019
rect 717 947 723 981
rect 757 947 763 981
rect 717 909 763 947
rect 717 875 723 909
rect 757 875 763 909
rect 717 837 763 875
rect 717 803 723 837
rect 757 803 763 837
rect 717 765 763 803
rect 717 731 723 765
rect 757 731 763 765
rect 717 693 763 731
rect 717 659 723 693
rect 757 659 763 693
rect 717 621 763 659
rect 717 587 723 621
rect 757 587 763 621
rect 717 549 763 587
rect 717 515 723 549
rect 757 515 763 549
rect 717 477 763 515
rect 717 443 723 477
rect 757 443 763 477
rect 717 405 763 443
rect 717 371 723 405
rect 757 371 763 405
rect 717 355 763 371
rect 1175 1629 1221 1645
rect 1175 1595 1181 1629
rect 1215 1595 1221 1629
rect 1175 1557 1221 1595
rect 1175 1523 1181 1557
rect 1215 1523 1221 1557
rect 1175 1485 1221 1523
rect 1175 1451 1181 1485
rect 1215 1451 1221 1485
rect 1175 1413 1221 1451
rect 1175 1379 1181 1413
rect 1215 1379 1221 1413
rect 1175 1341 1221 1379
rect 1175 1307 1181 1341
rect 1215 1307 1221 1341
rect 1175 1269 1221 1307
rect 1175 1235 1181 1269
rect 1215 1235 1221 1269
rect 1175 1197 1221 1235
rect 1175 1163 1181 1197
rect 1215 1163 1221 1197
rect 1175 1125 1221 1163
rect 1175 1091 1181 1125
rect 1215 1091 1221 1125
rect 1175 1053 1221 1091
rect 1175 1019 1181 1053
rect 1215 1019 1221 1053
rect 1175 981 1221 1019
rect 1175 947 1181 981
rect 1215 947 1221 981
rect 1175 909 1221 947
rect 1175 875 1181 909
rect 1215 875 1221 909
rect 1175 837 1221 875
rect 1175 803 1181 837
rect 1215 803 1221 837
rect 1175 765 1221 803
rect 1175 731 1181 765
rect 1215 731 1221 765
rect 1175 693 1221 731
rect 1175 659 1181 693
rect 1215 659 1221 693
rect 1175 621 1221 659
rect 1175 587 1181 621
rect 1215 587 1221 621
rect 1175 549 1221 587
rect 1175 515 1181 549
rect 1215 515 1221 549
rect 1175 477 1221 515
rect 1175 443 1181 477
rect 1215 443 1221 477
rect 1175 405 1221 443
rect 1175 371 1181 405
rect 1215 371 1221 405
rect 1175 355 1221 371
rect 1633 1629 1679 1645
rect 1633 1595 1639 1629
rect 1673 1595 1679 1629
rect 1633 1557 1679 1595
rect 1633 1523 1639 1557
rect 1673 1523 1679 1557
rect 1633 1485 1679 1523
rect 1633 1451 1639 1485
rect 1673 1451 1679 1485
rect 1633 1413 1679 1451
rect 1633 1379 1639 1413
rect 1673 1379 1679 1413
rect 1633 1341 1679 1379
rect 1633 1307 1639 1341
rect 1673 1307 1679 1341
rect 1633 1269 1679 1307
rect 1633 1235 1639 1269
rect 1673 1235 1679 1269
rect 1633 1197 1679 1235
rect 1633 1163 1639 1197
rect 1673 1163 1679 1197
rect 1633 1125 1679 1163
rect 1633 1091 1639 1125
rect 1673 1091 1679 1125
rect 1633 1053 1679 1091
rect 1633 1019 1639 1053
rect 1673 1019 1679 1053
rect 1633 981 1679 1019
rect 1633 947 1639 981
rect 1673 947 1679 981
rect 1633 909 1679 947
rect 1633 875 1639 909
rect 1673 875 1679 909
rect 1633 837 1679 875
rect 1633 803 1639 837
rect 1673 803 1679 837
rect 1633 765 1679 803
rect 1633 731 1639 765
rect 1673 731 1679 765
rect 1633 693 1679 731
rect 1633 659 1639 693
rect 1673 659 1679 693
rect 1633 621 1679 659
rect 1633 587 1639 621
rect 1673 587 1679 621
rect 1633 549 1679 587
rect 1633 515 1639 549
rect 1673 515 1679 549
rect 1633 477 1679 515
rect 1633 443 1639 477
rect 1673 443 1679 477
rect 1633 405 1679 443
rect 1633 371 1639 405
rect 1673 371 1679 405
rect 1633 355 1679 371
rect 2091 1629 2137 1645
rect 2091 1595 2097 1629
rect 2131 1595 2137 1629
rect 2091 1557 2137 1595
rect 2091 1523 2097 1557
rect 2131 1523 2137 1557
rect 2091 1485 2137 1523
rect 2091 1451 2097 1485
rect 2131 1451 2137 1485
rect 2091 1413 2137 1451
rect 2091 1379 2097 1413
rect 2131 1379 2137 1413
rect 2091 1341 2137 1379
rect 2091 1307 2097 1341
rect 2131 1307 2137 1341
rect 2091 1269 2137 1307
rect 2091 1235 2097 1269
rect 2131 1235 2137 1269
rect 2091 1197 2137 1235
rect 2091 1163 2097 1197
rect 2131 1163 2137 1197
rect 2091 1125 2137 1163
rect 2091 1091 2097 1125
rect 2131 1091 2137 1125
rect 2091 1053 2137 1091
rect 2091 1019 2097 1053
rect 2131 1019 2137 1053
rect 2091 981 2137 1019
rect 2091 947 2097 981
rect 2131 947 2137 981
rect 2091 909 2137 947
rect 2091 875 2097 909
rect 2131 875 2137 909
rect 2091 837 2137 875
rect 2091 803 2097 837
rect 2131 803 2137 837
rect 2091 765 2137 803
rect 2091 731 2097 765
rect 2131 731 2137 765
rect 2091 693 2137 731
rect 2091 659 2097 693
rect 2131 659 2137 693
rect 2091 621 2137 659
rect 2091 587 2097 621
rect 2131 587 2137 621
rect 2091 549 2137 587
rect 2091 515 2097 549
rect 2131 515 2137 549
rect 2091 477 2137 515
rect 2091 443 2097 477
rect 2131 443 2137 477
rect 2091 405 2137 443
rect 2091 371 2097 405
rect 2131 371 2137 405
rect 2091 355 2137 371
rect 2549 1629 2595 1645
rect 2549 1595 2555 1629
rect 2589 1595 2595 1629
rect 2549 1557 2595 1595
rect 2549 1523 2555 1557
rect 2589 1523 2595 1557
rect 2549 1485 2595 1523
rect 2549 1451 2555 1485
rect 2589 1451 2595 1485
rect 2549 1413 2595 1451
rect 2549 1379 2555 1413
rect 2589 1379 2595 1413
rect 2549 1341 2595 1379
rect 2549 1307 2555 1341
rect 2589 1307 2595 1341
rect 2549 1269 2595 1307
rect 2549 1235 2555 1269
rect 2589 1235 2595 1269
rect 2549 1197 2595 1235
rect 2549 1163 2555 1197
rect 2589 1163 2595 1197
rect 2549 1125 2595 1163
rect 2549 1091 2555 1125
rect 2589 1091 2595 1125
rect 2549 1053 2595 1091
rect 2549 1019 2555 1053
rect 2589 1019 2595 1053
rect 2549 981 2595 1019
rect 2549 947 2555 981
rect 2589 947 2595 981
rect 2549 909 2595 947
rect 2549 875 2555 909
rect 2589 875 2595 909
rect 2549 837 2595 875
rect 2549 803 2555 837
rect 2589 803 2595 837
rect 2549 765 2595 803
rect 2549 731 2555 765
rect 2589 731 2595 765
rect 2549 693 2595 731
rect 2549 659 2555 693
rect 2589 659 2595 693
rect 2549 621 2595 659
rect 2549 587 2555 621
rect 2589 587 2595 621
rect 2549 549 2595 587
rect 2549 515 2555 549
rect 2589 515 2595 549
rect 2549 477 2595 515
rect 2549 443 2555 477
rect 2589 443 2595 477
rect 2549 405 2595 443
rect 2549 371 2555 405
rect 2589 371 2595 405
rect 2549 355 2595 371
rect 3007 1629 3053 1645
rect 3007 1595 3013 1629
rect 3047 1595 3053 1629
rect 3007 1557 3053 1595
rect 3007 1523 3013 1557
rect 3047 1523 3053 1557
rect 3007 1485 3053 1523
rect 3007 1451 3013 1485
rect 3047 1451 3053 1485
rect 3007 1413 3053 1451
rect 3007 1379 3013 1413
rect 3047 1379 3053 1413
rect 3007 1341 3053 1379
rect 3007 1307 3013 1341
rect 3047 1307 3053 1341
rect 3007 1269 3053 1307
rect 3007 1235 3013 1269
rect 3047 1235 3053 1269
rect 3007 1197 3053 1235
rect 3007 1163 3013 1197
rect 3047 1163 3053 1197
rect 3007 1125 3053 1163
rect 3007 1091 3013 1125
rect 3047 1091 3053 1125
rect 3007 1053 3053 1091
rect 3007 1019 3013 1053
rect 3047 1019 3053 1053
rect 3007 981 3053 1019
rect 3007 947 3013 981
rect 3047 947 3053 981
rect 3007 909 3053 947
rect 3007 875 3013 909
rect 3047 875 3053 909
rect 3007 837 3053 875
rect 3007 803 3013 837
rect 3047 803 3053 837
rect 3007 765 3053 803
rect 3007 731 3013 765
rect 3047 731 3053 765
rect 3007 693 3053 731
rect 3007 659 3013 693
rect 3047 659 3053 693
rect 3007 621 3053 659
rect 3007 587 3013 621
rect 3047 587 3053 621
rect 3007 549 3053 587
rect 3007 515 3013 549
rect 3047 515 3053 549
rect 3007 477 3053 515
rect 3007 443 3013 477
rect 3047 443 3053 477
rect 3007 405 3053 443
rect 3007 371 3013 405
rect 3047 371 3053 405
rect 3007 355 3053 371
rect 120 17 3094 60
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3094 17
rect 120 -60 3094 -17
<< labels >>
flabel locali s 3034 104 3094 164 1 FreeSans 1250 0 0 0 GATE
port 1 nsew
flabel locali s 3034 1690 3094 1730 1 FreeSans 1250 0 0 0 SOURCE
port 2 nsew
flabel locali s 3034 210 3094 270 1 FreeSans 1250 0 0 0 DRAIN
port 3 nsew
flabel nwell s 120 1850 180 1910 1 FreeSans 1250 0 0 0 VPWR
port 4 nsew
flabel metal1 s 120 -30 278 30 1 FreeSans 1250 0 0 0 VGND
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 3395 1880
<< end >>
